/*****************************************************************************/
//
// Module          : cae_mc_rdord.vpp
// Revision        :  Revision: 1.12  
// Last Modified On:  Date: 2013-02-26 18:37:09  
// Last Modified By:  Author: gedwards  
//
//-----------------------------------------------------------------------------
//
// Original Author : gedwards
// Created On      : Wed Oct 10 09:26:08 2007
//
//-----------------------------------------------------------------------------
//
// Description     : Read ordering cache for MC loads
//
//-----------------------------------------------------------------------------
//
// Copyright (c) 2007 : created by Convey Computer Corp. This model is the
// confidential and proprietary property of Convey Computer Corp.
//
/*****************************************************************************/
/*  Id: cae_mc_rdord.vpp,v 1.12 2013-02-26 18:37:09 gedwards Exp   */

`timescale 1 ns / 1 ps

(* keep_hierarchy = "true" *)
module cae_mc_rdord (/*AUTOARG*/
   // Outputs
   p_rq_stall, m_rq_bus, m_rq_vld, m_rq_flush, m_rs_stall, p_rs_vld,
   p_rs_bus, p_rs_flush_cmplt,
   // Inputs
   clk2x, clk, i_reset, p_rq_bus, p_rq_vld, p_rq_flush, m_rq_stall,
   m_rs_vld, m_rs_bus, m_rs_flush_cmplt, p_rs_stall
   ) ;
  
   /* ----------         include files        ---------- */
  // Generated by src/generate_ae_fpxbar.pl in efox/project_bfms/Ae_FpXbar
/*****************************************************************************/
//
// Module     : aemc_messages.vh
// Revision   :  Revision: 1.11  
//
//-----------------------------------------------------------------------------
//
// Description: Convey ae_mc message encodings - EFox Project
//
//-----------------------------------------------------------------------------
//
// Copyright (c) 2007-2012 by Convey Computer Corp. This file is
// the confidential and proprietary property of Convey Computer Corp.
//
/*****************************************************************************/
//  Id: aemc_messages.vh,v 1.11 2014/05/22 21:09:06 gedwards Exp  

// AeMc AE_Rq format
`define AE_RQ_CMD               2:0
`define AE_RQ_RSVD1             5:3
`define AE_RQ_TID              15:6
`define AE_RQ_SUB             19:16
`define AE_RQ_RSVD0           21:20
`define AE_RQ_LEN             23:22
`define AE_RQ_VADR            71:24

// AeMc AE_Data format
`define AE_DATA_CMD             2:0
`define AE_DATA_RSVD1           5:3
`define AE_DATA_RSVD0           7:6
`define AE_DATA_DATA           71:8

// AeMc AE_Mc_null format
`define AE_MC_NULL_CMD          2:0

// McAe MC_Ae_null format
`define MC_AE_NULL_CMD          2:0

// McAe AE_Rs format
`define AE_RS_CMD               2:0
`define AE_RS_SUB               5:3
`define AE_RS_TID              15:6
`define AE_RS_DATA            79:16

// PDK AE_Rq format
`define PDK_RQ_CMD               2:0
`define PDK_RQ_SUB               6:3
`define PDK_RQ_LEN               8:7
`define PDK_RQ_VADR             56:9
`define PDK_RQ_DATA           120:57
`define PDK_RQ_RTNCTL        152:121
`define PDK_RQ_MSB_LSB         152:0

// PDK AE_Rs format
`define PDK_RS_CMD               2:0
`define PDK_RS_SUB               5:3 //rs_sub = rq_sub[3:1], for IFETCH it has vadr[5:3]
`define PDK_RS_DATA             69:6
`define PDK_RS_RTNCTL         101:70
`define PDK_RS_MSB_LSB         101:0

localparam
	// AEMC command types
	AEMC_CMD_IDLE         = 3'd0,
	AEMC_CMD_RD           = 3'd1,
	AEMC_CMD_WR           = 3'd2,
	AEMC_CMD_FENCE        = 3'd3,
	AEMC_CMD_FE           = 3'd4,
	AEMC_CMD_ATOMIC       = 3'd5,
	AEMC_CMD_RESERVED     = 3'd6,
	AEMC_CMD_IFETCH       = 3'd7,

	// Names used for HC and WX
        AEMC_CMD_RD8            = 3'd1,
        AEMC_CMD_WR8            = 3'd2,
        AEMC_CMD_WR64           = 3'd6,
        AEMC_CMD_RD64           = 3'd7,

	// AEMC Rd - sub cmd
	AEMC_CMD_RD_BYTE      = 4'd0,

	// AEMC Wr - sub cmd
	AEMC_CMD_WR_BYTE      = 4'd0,
	AEMC_CMD_WR_64_BYTE   = 4'd1,

	// AEMC FE - sub cmd
	AEMC_CMD_FE_RFE       = 4'd0,
	AEMC_CMD_FE_RFF       = 4'd1,
	AEMC_CMD_FE_FAD       = 4'd2,
	AEMC_CMD_FE_REF       = 4'd3,
	AEMC_CMD_FE_WEF       = 4'd4,
	AEMC_CMD_FE_WFF       = 4'd5,
	AEMC_CMD_FE_WXF       = 4'd6,
	AEMC_CMD_FE_WXE       = 4'd7,
	AEMC_CMD_FE_RXX       = 4'd8,
	AEMC_CMD_FE_PUR       = 4'd12,

	// AEMC Atomic - sub cmd
	AEMC_CMD_ATOM_ADD     = 4'd0,
	AEMC_CMD_ATOM_SUB     = 4'd1,
	AEMC_CMD_ATOM_EXCH    = 4'd2,
	AEMC_CMD_ATOM_MIN     = 4'd3,
	AEMC_CMD_ATOM_MAX     = 4'd4,
	AEMC_CMD_ATOM_INC     = 4'd5,
	AEMC_CMD_ATOM_DEC     = 4'd6,
	AEMC_CMD_ATOM_AND     = 4'd7,
	AEMC_CMD_ATOM_OR      = 4'd8,
	AEMC_CMD_ATOM_XOR     = 4'd9,
	AEMC_CMD_ATOM_CAS     = 4'd10,

	// MCAE command types
	MCAE_CMD_IDLE         = 3'd0,
	MCAE_CMD_RD_DATA      = 3'd2,
	MCAE_CMD_WR_CMP       = 3'd3,  // WR8 complete for Fox
	MCAE_CMD_FE_RETRY     = 3'd4,
	MCAE_CMD_FE_DATA      = 3'd5,
	MCAE_CMD_ATOMIC_DATA  = 3'd6,
	MCAE_CMD_IFILL        = 3'd7,

        // New names for HC and WX
        MCAE_CMD_WR64_CMP     = 3'd1,   // placeholder for Fox platform
        MCAE_CMD_RD8_DATA     = 3'd2,
        MCAE_CMD_RD64_DATA    = 3'd7,

	// ae size field
	MC_SIZE_BYTE          = 2'd0,
	MC_SIZE_WORD          = 2'd1,
	MC_SIZE_LONG          = 2'd2,
	MC_SIZE_QUAD          = 2'd3;



   parameter MC_READ_ORDER = 0;
   parameter MC_WR_CMP_IF = 0;
   parameter RDCTL_TOP = 23;
   parameter RDCTL_BITS = 10;
   parameter RDCTL_BOTTOM = RDCTL_TOP-RDCTL_BITS+1;

   /* ----------        port declarations     ---------- */

    input		clk2x;
    input		clk;
    input		i_reset;

    // REQUEST FLOW ======================
    // Personality-side interface ----
    input [`PDK_RQ_MSB_LSB] p_rq_bus;
    input		                p_rq_vld;
    input		                p_rq_flush;
    output		              p_rq_stall;

    // MC/XB-side interface --------
    output [`PDK_RQ_MSB_LSB] m_rq_bus;
    output		               m_rq_vld;
    output		               m_rq_flush;
    input		               m_rq_stall;
   
    // RESPONSE FLOW ======================
    // MC/XB-side interface --------
    input		                m_rs_vld;
    input [`PDK_RS_MSB_LSB] m_rs_bus;
    output		              m_rs_stall;
    input		                m_rs_flush_cmplt; 

    // Personality-side interface ----
    //
    output		               p_rs_vld;
    output [`PDK_RS_MSB_LSB] p_rs_bus;
    input		                 p_rs_stall;
    output		               p_rs_flush_cmplt;
//   output		csr_txns_out;
//   output		csr_txns_hld;

   /* ----------          wires & regs        ---------- */

   wire		      reset;
   reg          r_t1_rq_vld;
   reg  [1:0]   r_t1_rq_len;
   reg  [2:0]   r_t1_rq_cmd;
   reg  [3:0]   r_t1_rq_sub;
   reg  [47:0]  r_t1_rq_vadr;
   reg  [63:0]  r_t1_rq_data;
   reg  [31:0]  r_t1_rq_rtnctl;
   reg  [31:0]  c_t1_rq_rtnctl;
   reg          r_t1_rq_flush;
   reg          r_t2_rq_vld;
   reg  [1:0]   r_t2_rq_len;
   reg  [2:0]   r_t2_rq_cmd;
   reg  [3:0]   r_t2_rq_sub;
   reg  [47:0]  r_t2_rq_vadr;
   reg  [63:0]  r_t2_rq_data;
   reg  [31:0]  r_t2_rq_rtnctl;
   reg          r_t2_rq_flush;

   wire  [8:0]   c_t0_rq_tid;
   reg   [8:0]   r_t1_rq_tid;
   reg   [8:0]   r_t2_rq_tid;
   reg   [8:0]   r_t3_rq_tid;

   wire  [8:0]   c_t0_rptr;
	(* shreg_extract = "no" *)
	(* equivalent_register_removal = "no" *)
	(* S = "TRUE" *)
	(* KEEP = "TRUE" *)
   reg   [8:0]   r_t1_rptr, r_t1_rptr1;
   reg   [9:0]   c_tid_free_cnt;
   reg   [9:0]   r_tid_free_cnt;
   reg   [9:0]   c_txns_out_cnt;
   reg   [9:0]   r_txns_out_cnt;

    reg	 r_p_rs_stall;

    wire c_t1_dout_vld;

    wire [76:0]	bram_dout;
    wire [3:0]	fifo_cnt;
    wire		fifo_full;
    wire		fifo_empty;
    wire		fifo_push;
    reg 		r_fifo_push;
    wire		c_t1_ram_toggle;
    reg 		r_t1_ram_toggle;

    reg pend_ram [511:0];
    reg recd_ram [511:0];

    wire rd_pending;
    wire rd_returned;
    wire c_t1_pend_we;
    wire c_t1_recd_we;

    wire          c_p_rs_vld;
    reg           r_p_rs_vld;
    wire [2:0]    c_p_rs_cmd;
    reg  [2:0]    r_p_rs_cmd;
    wire [2:0]    c_p_rs_sub;
    reg  [2:0]    r_p_rs_sub;
    wire [6:0]    c_p_rs_rtnctl;
    reg  [6:0]    r_p_rs_rtnctl;
    wire [63:0]	  c_p_rs_data;
    reg  [63:0]	  r_p_rs_data;
    
    // Signal breakout for debussy/ possibly for code...
    wire [2:0]  p_rq_cmd    = p_rq_bus[`PDK_RQ_CMD];
    wire [3:0]  p_rq_sub    = p_rq_bus[`PDK_RQ_SUB];
    wire [1:0]  p_rq_len    = p_rq_bus[`PDK_RQ_LEN];
    wire [47:0] p_rq_vadr   = p_rq_bus[`PDK_RQ_VADR];
    wire [63:0] p_rq_data   = p_rq_bus[`PDK_RQ_DATA];
    wire [31:0] p_rq_rtnctl = p_rq_bus[`PDK_RQ_RTNCTL];
    // Response decode
    wire [2:0]  m_rs_cmd    = m_rs_bus[`PDK_RS_CMD];
    wire [3:0]  m_rs_sub    = m_rs_bus[`PDK_RS_SUB];
    wire [63:0] m_rs_data   = m_rs_bus[`PDK_RS_DATA];
    wire [31:0] m_rs_rtnctl = m_rs_bus[`PDK_RS_RTNCTL];
    wire m_rs_ld = (m_rs_cmd==MCAE_CMD_RD_DATA)&&m_rs_vld;
    wire m_rs_st = (m_rs_cmd==MCAE_CMD_WR_CMP)&&m_rs_vld;
   /* ----------      combinatorial blocks    ---------- */

generate if (MC_READ_ORDER == 0) begin : gno_rdord
    assign m_rq_bus = p_rq_bus;
    assign m_rq_vld = p_rq_vld;
    assign m_rq_flush = p_rq_flush;
    assign p_rq_stall = m_rq_stall;
    assign m_rs_stall = p_rs_stall;
    assign p_rs_vld = m_rs_vld;
    assign p_rs_bus = m_rs_bus;
    assign p_rs_flush_cmplt = m_rs_flush_cmplt;
//   assign csr_txns_out = 1'b0;
//   assign csr_txns_hld = 1'b0;
end else begin : grdord
    // wire/regs only for rd-order case 
    wire        c_p_rq_stall;
    reg         r_p_rq_stall;
    wire  [8:0] c_t1_pend_wptr;
    wire  [8:0] c_t1_recd_wptr;
    wire  [8:0] c_rst_cnt;
    reg   [8:0] r_rst_cnt;
    reg         r_t2_recd_we;
    wire        c_t2_recd_we;
    reg  [8:0]  r_t2_recd_wptr;
    reg         r_t2_rs_ramtoggle;

    // response path
    reg		r_t1_rs_vld;
    reg  [31:0] r_t1_rs_rtnctl;
    reg  [63:0] r_t1_rs_data;
    reg  [2:0]  r_t1_rs_cmd;
    reg  [2:0]  r_t1_rs_sub;
    reg         r_cutoff;

    // output port assignments    
    // RQ flow
    assign m_rq_vld = r_t2_rq_vld;
    assign m_rq_bus[`PDK_RQ_CMD]    = r_t2_rq_cmd;
    assign m_rq_bus[`PDK_RQ_SUB]    = r_t2_rq_sub;
    assign m_rq_bus[`PDK_RQ_LEN]    = r_t2_rq_len;
    assign m_rq_bus[`PDK_RQ_VADR]   = r_t2_rq_vadr;
    assign m_rq_bus[`PDK_RQ_DATA]   = r_t2_rq_data;
    assign m_rq_bus[`PDK_RQ_RTNCTL] = r_t2_rq_rtnctl;
    assign m_rq_flush = r_t2_rq_flush;
    assign p_rq_stall = r_p_rq_stall;
    // RS flow
    assign p_rs_bus[`PDK_RS_CMD] = r_p_rs_cmd;
    assign p_rs_bus[`PDK_RS_SUB] = r_p_rs_sub;
    assign p_rs_bus[`PDK_RS_DATA] = r_p_rs_data;
    assign p_rs_bus[`PDK_RS_RTNCTL] = {25'b0,r_p_rs_rtnctl};
    
if (MC_WR_CMP_IF == 0) begin : gflush
    // With the flush interface invoked, no point in sending the wr-rsp's back 
    // throught the async block, so squash them here
    assign p_rs_vld = r_p_rs_vld && (r_p_rs_cmd==MCAE_CMD_RD_DATA);
end else begin : gwrcmp 
    // need to return wr_cmps to the personality
    assign p_rs_vld = r_p_rs_vld;
end
    
    assign m_rs_stall = 1'b0;
    reg r_m_rs_flush_cmplt;
    always @(posedge clk2x) begin
      r_m_rs_flush_cmplt <= m_rs_flush_cmplt;
    end
    assign p_rs_flush_cmplt = r_m_rs_flush_cmplt;

    // Set certain rtnctl bits to track where we stored this request in the
    // ordering RAMs
    always @* begin
      c_t1_rq_rtnctl = r_t1_rq_rtnctl;
      if (r_t1_rq_vld)
        c_t1_rq_rtnctl[RDCTL_TOP:RDCTL_BOTTOM] = {r_t1_ram_toggle,r_t1_rq_tid};
    end

    // RQ Stall logic ---------- 
    // If we are stalled by xb/mc or our tid_free_cnt is <9, stall personality
    assign c_p_rq_stall = m_rq_stall || (r_tid_free_cnt < 'd9);

    // logic to determine when to shutoff pulling pushing responses from DRAMS
    // into rsp fifos
    wire c_cutoff = (r_txns_out_cnt <= 'd0) ||
                    ((r_txns_out_cnt == 'd1) && r_fifo_push); 
  
    assign c_t1_dout_vld =  (rd_pending==rd_returned) && ~c_cutoff;
    assign fifo_push = c_t1_dout_vld && (fifo_cnt < 4'd4);

    assign c_t1_pend_we = r_t1_rq_vld | reset;

    assign c_t1_pend_wptr = reset ? r_rst_cnt : r_t1_rq_tid;
    assign c_t1_recd_wptr = reset ? r_rst_cnt : r_t1_rs_rtnctl[RDCTL_TOP-1:RDCTL_BOTTOM];
    // leda W484 off
    assign c_rst_cnt = r_rst_cnt + 'd1;
    // leda W484 on

    assign c_t1_ram_toggle = (r_t1_rq_tid == 'd511) && r_t1_rq_vld ? ~r_t1_ram_toggle : r_t1_ram_toggle;

    always @(posedge clk2x) begin
      if (c_t1_pend_we)
        pend_ram[c_t1_pend_wptr] <= reset | r_t1_ram_toggle;
    end

    // RS pipe ----------------
    assign c_t1_recd_we = r_t1_rs_vld; // currently order both RD&WR
    assign c_t2_recd_we = r_t2_recd_we | reset;

    always @(posedge clk2x) begin
      if (c_t2_recd_we)
        recd_ram[r_t2_recd_wptr] <= reset | r_t2_rs_ramtoggle;
    end

    assign rd_pending = pend_ram[r_t1_rptr1];
    assign rd_returned = recd_ram[r_t1_rptr1];

    // leda W484 off
    always @* begin
      // r_p_rs_vld includes ALL responses ... fixme if changing to RDONLY
      // ordering
      case ({r_t1_rq_vld, r_p_rs_vld})
      2'b00:  c_tid_free_cnt = r_tid_free_cnt;
      2'b01:  c_tid_free_cnt = r_tid_free_cnt + 'b1;
      2'b10:  c_tid_free_cnt = r_tid_free_cnt - 'b1;
      2'b11:  c_tid_free_cnt = r_tid_free_cnt;
      endcase
   end
   
    always @* begin
      case ({r_t2_rq_vld, r_fifo_push})
      2'b00:  c_txns_out_cnt = r_txns_out_cnt;
      2'b01:  c_txns_out_cnt = r_txns_out_cnt - 'b1;
      2'b10:  c_txns_out_cnt = r_txns_out_cnt + 'b1;
      2'b11:  c_txns_out_cnt = r_txns_out_cnt;
      endcase
    end

   //assign c_t0_rptr = r_t1_rptr + {8'b0,fifo_push};
   assign c_t0_rptr = r_t1_rptr + 'b1;
   assign c_t0_rq_tid = r_t1_rq_tid + 'b1;
  // leda W484 on

   sdpram #(.DEPTH(512),.WIDTH(3+3+7+64),.PIPE(0)) dpram (
      .clk      (clk2x),
      .din      ({r_t1_rs_sub[2:0], r_t1_rs_cmd[2:0],r_t1_rs_rtnctl[6:0], r_t1_rs_data[63:0]}),
      .wadr     (c_t1_recd_wptr),
      .we       (c_t1_recd_we),
      .radr     (r_t1_rptr),
      .ce       (1'b1),
      .oreg_ce  (1'b1),
      .oreg_rst (1'b0),
      .dout     (bram_dout[76:0])
   );

   assign c_p_rs_vld = !fifo_empty && !r_p_rs_stall;

  // leda B_1011 off
   fifo #(.DEPTH(8), .WIDTH(3+3+7+64)) rsp_fifo (
    .clk    (clk2x),
    .reset  (reset),
    .push   (r_fifo_push),
    .din    (bram_dout),
    .afull  (),
    .full   (fifo_full),
    .cnt    (fifo_cnt),
    .oclk   (clk2x),
    .pop    (c_p_rs_vld),
    .dout   ({c_p_rs_sub[2:0], c_p_rs_cmd[2:0], c_p_rs_rtnctl[6:0], c_p_rs_data[63:0]}),
    .empty  (fifo_empty),
    .rcnt   ()
   );
  // leda B_1011 on

   // debug 
/*
   wire  [63:0]  c_out_cnt, r_out_cnt;
   wire  [63:0]  c_hld_cnt, r_hld_cnt;
   wire c_txns_out, r_txns_out;
   wire c_txns_hld, r_txns_hld;

   assign c_out_cnt = r_out_cnt + r_t1_rq_vld - r_t1_rs_vld;
   assign c_hld_cnt = r_hld_cnt + r_t1_rs_vld - p_rs_vld;

   assign c_txns_out = r_out_cnt > 'd0;
   assign c_txns_hld = r_hld_cnt > 'd0;

   DFFC(64, reg_out_cnt, clk2x, reset, c_out_cnt, r_out_cnt);
   DFFC(64, reg_hld_cnt, clk2x, reset, c_hld_cnt, r_hld_cnt);
   DFF ( 1, reg_txns_out, clk2x, c_txns_out, r_txns_out);
   DFF ( 1, reg_txns_hld, clk2x, c_txns_hld, r_txns_hld);
   DFF ( 1, reg_csr_txns_out, clk_csr, r_txns_out, csr_txns_out);
   DFF ( 1, reg_csr_txns_hld, clk_csr, r_txns_hld, csr_txns_hld);
*/
   /* ----------      external module calls   ---------- */


  /* ----------            registers         ---------- */

  // register request from personality
  always @(posedge clk2x) begin
    r_t2_recd_we <= c_t1_recd_we;
    r_t2_recd_wptr <= c_t1_recd_wptr;
    r_t2_rs_ramtoggle <= r_t1_rs_rtnctl[RDCTL_TOP];
   
    r_cutoff <= reset ? 1'b1 : c_cutoff;
    r_fifo_push <= reset ? 1'b0 : fifo_push;

    r_p_rq_stall <= reset ? 1'b0 : c_p_rq_stall;

    r_t1_rq_vld <= reset ? 1'b0 : p_rq_vld;
    r_t1_rq_len <= reset ? 2'b0 : p_rq_len;
    r_t1_rq_cmd <= reset ? 3'b0 : p_rq_cmd;
    r_t1_rq_sub <= reset ? 4'b0 : p_rq_sub;
    r_t1_rq_vadr <= reset ? 48'b0 : p_rq_vadr;
    r_t1_rq_data <= reset ? 64'b0 : p_rq_data;
    r_t1_rq_rtnctl <= reset ? 32'b0 : p_rq_rtnctl;
    r_t1_rq_flush <= reset ? 1'b0 : p_rq_flush;

    // second rq-pipe stage    
    r_t2_rq_vld <= reset ? 1'b0 : r_t1_rq_vld;
    r_t2_rq_len <= reset ? 2'b0 : r_t1_rq_len;
    r_t2_rq_cmd <= reset ? 3'b0 : r_t1_rq_cmd;
    r_t2_rq_sub <= reset ? 4'b0 : r_t1_rq_sub;
    r_t2_rq_vadr <= reset ? 48'b0 : r_t1_rq_vadr;
    r_t2_rq_data <= reset ? 64'b0 : r_t1_rq_data;
    r_t2_rq_rtnctl <= reset ? 32'b0 : c_t1_rq_rtnctl;
    r_t2_rq_flush <= reset ? 1'b0 : r_t1_rq_flush;

    // grab the incremented rq-tid whenever we see a new rq-load
    r_t1_rq_tid <= reset ? 'b0 : r_t1_rq_vld ? c_t0_rq_tid : r_t1_rq_tid;
    r_t2_rq_tid <= reset ? 'b0 : r_t1_rq_tid;
    r_t3_rq_tid <= reset ? 'b0 : r_t2_rq_tid;
   
    r_t1_ram_toggle <= reset ? 1'b0 : c_t1_ram_toggle;

    // response pipe
    r_t1_rs_vld <= reset ? 1'b0 : m_rs_vld;
    r_t1_rs_rtnctl <= reset ? 32'b0 : m_rs_rtnctl;
    r_t1_rs_data <= reset ? 64'b0 : m_rs_data;
    r_t1_rs_cmd <= reset ? 3'b0 : m_rs_cmd;
    r_t1_rs_sub <= reset ? 3'b0 : m_rs_sub;
    
    // response pipe, from rs-fifo to rs-outputs
    r_p_rs_rtnctl <= c_p_rs_rtnctl;
    r_p_rs_cmd <= c_p_rs_cmd;
    r_p_rs_sub <= c_p_rs_sub;
    r_p_rs_data <= c_p_rs_data; 

    // rs stall
    r_p_rs_stall <= p_rs_stall;   
    r_p_rs_vld <= c_p_rs_vld;
   
    r_rst_cnt <= c_rst_cnt;
  
    r_tid_free_cnt <= reset ? 'd512 : c_tid_free_cnt;
    r_txns_out_cnt <= reset ? 'b0   : c_txns_out_cnt; 
   
    //r_t1_rptr <= reset ? 9'b0 : c_t0_rptr;
    r_t1_rptr <= reset ? 'b0 : fifo_push ? c_t0_rptr : r_t1_rptr;
    r_t1_rptr1 <= reset ? 'b0 : fifo_push ? c_t0_rptr : r_t1_rptr1;
  end
   reset_flop_1 reg_reset ( .clk(clk), .i_reset(i_reset), .reset(reset) );

   // synopsys translate_off

   // Parameters: 1-Severity: Don't Stop, 2-start check only after negedge of reset
   assert_never #(0, 2, "***ERROR ASSERT:  Read Order TID underflow") 
     a0 (.clk(clk2x), .reset_n(~reset), .test_expr((r_tid_free_cnt == 'd0) && r_t1_rq_vld));

   assert_never #(0, 2, "***ERROR ASSERT:  Read Order TID overflow") 
     a1 (.clk(clk2x), .reset_n(~reset), .test_expr((r_tid_free_cnt == 'd512) && r_p_rs_vld));

    // synopsys translate_on
end
endgenerate

endmodule // cae_mc_rdord

// This is the search path for the autoinst commands in emacs.
// After modification you must save file, then reld with C-x C-v
//
// Local Variables:
// verilog-library-directories:("." "../../common/xilinx") 
// verilog-library-flags:("-y ../../../REVISIONS/MX/common/lib -y ../../../REVISIONS/MX/common/xilinx -y ../../../REVISIONS/MX/project_common/lib")
// End:

